library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity decoder_5to32 is
Port ( a : in  STD_LOGIC_VECTOR (4 downto 0);
           y : out  STD_LOGIC_VECTOR (31 downto 0));
end decoder_5to32;

architecture Behavioral of decoder_5to32 is

begin
 process(a)
  begin
    case a is
		when "00000" =>
			y <= "00000000000000000000000000000001";
      when "00001" =>
        y <= "00000000000000000000000000000010";
		when "00010" =>
        y <= "00000000000000000000000000000100";
		when "00011" =>
        y <= "00000000000000000000000000001000";
      when "00100" =>
        y <= "00000000000000000000000000010000";
      when "00101" =>
        y <= "00000000000000000000000000100000";
		 when "00110" =>
		y <= "00000000000000000000000001000000";
		when "00111" =>
        y <= "00000000000000000000000010000000";
      when "01000" =>
        y <= "00000000000000000000000100000000";
      when "01001" =>
        y <= "00000000000000000000001000000000";
      when "01010" =>
        y <= "00000000000000000000010000000000";
		 when "01011" =>
		 y <= "00000000000000000000100000000000";
      when "01100" =>
        y <= "00000000000000000001000000000000";
		when "01101" =>
        y <= "00000000000000000010000000000000";
      when "01110" =>
        y <= "00000000000000000100000000000000";
      when "01111" =>
        y <= "00000000000000001000000000000000";  
		when "10000" =>
        y <= "00000000000000010000000000000000";
      when "10001" =>
        y <= "00000000000000100000000000000000";
      when "10010" =>
		 y <= "00000000000001000000000000000000";
		when "10011" =>
        y <= "00000000000010000000000000000000";
      when "10100" =>
        y <= "00000000000100000000000000000000";
      when "10101" =>
        y <= "00000000001000000000000000000000";
      when "10110" =>
        y <= "00000000010000000000000000000000";
      when "10111" =>
        y <= "00000000100000000000000000000000";
		when "11000" =>
			 y <= "00000001000000000000000000000000";
		  when "11001" =>
			 y <= "00000010000000000000000000000000";
		  when "11010" =>
			 y <= "00000100000000000000000000000000";
		  when "11011" =>
			 y <= "00001000000000000000000000000000";
		  when "11100" =>
			 y <= "00010000000000000000000000000000";
		  when "11101" =>
			 y <= "00100000000000000000000000000000";
		  when "11110" =>
			 y <= "01000000000000000000000000000000";
		  when "11111" =>
			 y <= "10000000000000000000000000000000"; 
		  when others =>
			y <=	"00000000000000000000000000000000";
		end case;
	end process;

end Behavioral;

